 constant scp  : std_logic_vector(31 downto 0) := (x"00000101");
 constant scp2 : std_logic_vector(31 downto 0) := (x"00000102");
 constant scp3 : std_logic_vector(31 downto 0) := (x"00000103");
 constant scp4 : std_logic_vector(31 downto 0) := (x"00000104");
 constant scp5 : std_logic_vector(31 downto 0) := (x"00000105");
 constant scp6 : std_logic_vector(31 downto 0) := (x"00000106");
 constant scp7 : std_logic_vector(31 downto 0) := (x"00000107");
 constant scp8 : std_logic_vector(31 downto 0) := (x"00000108");
 constant scp9 : std_logic_vector(31 downto 0) := (x"00000109");
     when scp => 
          mem_addr <= sp-1; sp <= sp-1;--init pop source address
                we <= "0"; -- enable read next state
        ir <= scp2;
          when scp2 => -- mem_addr updated
          mem_addr <= sp-1; sp <= sp-1;--init pop dest address
        we <= "0"; -- read
        ir <= scp3; -- one additional latency when simulate
              --ir <= scp4; -- HW ip skip sl3 
          when scp3 => -- douta not valid latency 1
                we <= "0"; -- read
                ir <= scp4;            
          when scp4 => -- douta valid
        we <= "0"; -- read
        ir <= scp5;     
          when scp5 => -- mem_data_out valid sourcxe addr
      mem_addr <= mem_data_out(A-1 downto 0);--source Address
        we <= "0"; -- read
                ir <= scp6;
          when scp6 => -- mem_addr updated, mem_data_out valid dest addr
        we <= "0"; -- read
        temp1 <= mem_data_out(A-1 downto 0);-- dest Address
        ir <= scp7; -- one additional latency when simulate
--              ir <= scp8; -- HW ip skip sl7
          when scp7 => -- douta not valid latency 1, 
                we <= "0"; -- read
                ir <= scp8;                    
          when scp8 => -- douta valid
        we <= "0"; -- read
        ir <= scp9;          
          when scp9 => -- mem_data_out valid
          mem_addr <= temp1; -- temp1 is dest addr
       mem_data_in <= mem_data_out;--source data
        we <= "1"; -- write enable in next state
               n_s <= fetch;
